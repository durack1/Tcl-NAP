netcdf geog {
dimensions:
	time = UNLIMITED ; // (24 currently)
	latitude = 59 ;
	longitude = 67 ;
variables:
	float time(time) ;
		time:_FillValue = nanf ;
		time:units = "days since 1700-1-1 0:0:0" ;
	float latitude(latitude) ;
		latitude:_FillValue = nanf ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:_FillValue = nanf ;
		longitude:units = "degrees_east" ;
	float tscrn(time, latitude, longitude) ;
		tscrn:_FillValue = nanf ;
		tscrn:long_name = "screen level (1.8m) temperature" ;
		tscrn:units = "K" ;
data:

 time = 95328, 95359, 95387, 95418, 95448, 95479, 95509, 95540, 95571, 95601, 
    95632, 95662, 95693, 95724, 95752, 95783, 95813, 95844, 95874, 95905, 
    95936, 95966, 95997, 96027 ;

 latitude = -48, -47.5, -47, -46.5, -46, -45.5, -45, -44.5, -44, -43.5, -43, 
    -42.5, -42, -41.5, -41, -40.5, -40, -39.5, -39, -38.5, -38, -37.5, -37, 
    -36.5, -36, -35.5, -35, -34.5, -34, -33.5, -33, -32.5, -32, -31.5, -31, 
    -30.5, -30, -29.5, -29, -28.5, -28, -27.5, -27, -26.5, -26, -25.5, -25, 
    -24.5, -24, -23.5, -23, -22.5, -22, -21.5, -21, -20.5, -20, -19.5, -19 ;

 longitude = 127, 127.5, 128, 128.5, 129, 129.5, 130, 130.5, 131, 131.5, 132, 
    132.5, 133, 133.5, 134, 134.5, 135, 135.5, 136, 136.5, 137, 137.5, 138, 
    138.5, 139, 139.5, 140, 140.5, 141, 141.5, 142, 142.5, 143, 143.5, 144, 
    144.5, 145, 145.5, 146, 146.5, 147, 147.5, 148, 148.5, 149, 149.5, 150, 
    150.5, 151, 151.5, 152, 152.5, 153, 153.5, 154, 154.5, 155, 155.5, 156, 
    156.5, 157, 157.5, 158, 158.5, 159, 159.5, 160 ;
}
