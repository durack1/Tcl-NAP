netcdf darlam {
dimensions:
	time = 24 ;
	y = 50 ;
	x = 44 ;
variables:
	float time(time) ;
		time:units = "days since 1700-1-1 0:0:0" ;
	float y(y) ;
	float x(x) ;
	float tscrn(time, y, x) ;
		tscrn:_FillValue = nanf ;
		tscrn:long_name = "screen level (1.8m) temperature" ;
		tscrn:units = "K" ;
data:

 time = 95328, 95359, 95387, 95418, 95448, 95479, 95509, 95540, 95571, 95601, 
    95632, 95662, 95693, 95724, 95752, 95783, 95813, 95844, 95874, 95905, 
    95936, 95966, 95997, 96027 ;

 y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 
    39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 
    39, 40, 41, 42, 43, 44 ;
}
