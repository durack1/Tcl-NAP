netcdf u {
dimensions:
	time = UNLIMITED ;
variables:
	float time(time) ;
data:
 time = 2, 4;
}
