netcdf lat_lon_60km {
dimensions:
	y = 50 ;
	x = 44 ;
variables:
	float latitude(y, x) ;
		latitude:units = "degrees_north" ;
	float longitude(y, x) ;
		longitude:units = "degrees_east" ;
	int x(x) ;
		x:_FillValue = -2147483648 ;
	int y(y) ;
		y:_FillValue = -2147483648 ;

// global attributes:
		:history = "25Feb2002 1245; bat064; text2nc lat_lon_60km.nc longitude\n",
    "25Feb2002 1245; bat064; text2nc lat_lon_60km.nc latitude\n",
    "" ;
data:

 x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 
    39, 40, 41, 42, 43, 44 ;

 y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 
    21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 
    39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;
}
